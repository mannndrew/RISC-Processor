module decoder
(

);

endmodule
