module SingleCycle;

endmodule