module regfile
(
	input write_data;
	input [4:0] read_address
	output read_data;
);